`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.10.2016 13:28:25
// Design Name: 
// Module Name: font_pong
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module word_pong(
    input [4:0] drom_addr_num,
    output reg [0:127] drom_data_num
);

always @(*)
    begin
	    case (drom_addr_num)
            0:drom_data_num = 128'b01111111111111111111111111110000000011111111111111111111111100000000111111111111111111111111000000001111111111111111111111111110;
            1:drom_data_num = 128'b01000000000000000000000000001000000100000000000000000000000010000001000000000000000000000000100000010000000000000000000000000000;
            2:drom_data_num = 128'b01000000000000000000000000000100001000000000000000000000000001000010000000000000000000000000010000100000000000000000000000000000;
            3:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
            4:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
            5:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
            6:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
            7:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
            8:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
            9:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
           10:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
           11:drom_data_num = 128'b01000000000000000000000000000010010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
           12:drom_data_num = 128'b01000000000000000000000000000100010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
           13:drom_data_num = 128'b01000000000000000000000000001000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000000;
           14:drom_data_num = 128'b01011111111111111111111111110000010000000000000000000000000000100100000000000000000000000000001001000011111111111111111111110000;
           15:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000001000;
           16:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000100;
           17:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           18:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           19:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           20:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           21:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           22:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           23:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           24:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           25:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           26:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           27:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           28:drom_data_num = 128'b01000000000000000000000000000000010000000000000000000000000000100100000000000000000000000000001001000000000000000000000000000010;
           29:drom_data_num = 128'b01000000000000000000000000000000001000000000000000000000000001000100000000000000000000000000001000100000000000000000000000000100;
           30:drom_data_num = 128'b01000000000000000000000000000000000100000000000000000000000010000100000000000000000000000000001000010000000000000000000000001000;
           31:drom_data_num = 128'b01000000000000000000000000000000000011111111111111111111111100000100000000000000000000000000001000001111111111111111111111110000;
        endcase
    end

endmodule