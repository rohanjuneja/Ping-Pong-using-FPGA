`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/19/2016 06:24:17 PM
// Design Name: 
// Module Name: font_number
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module font_ball(
    input [4:0] drom_addr_num,
    output reg [0:31] drom_data_num
);
    
always @(*) begin
        case (drom_addr_num)
            0:drom_data_num = 32'b00000000000000000000000000000000;
            1:drom_data_num = 32'b00000000000001111110000000000000;
            2:drom_data_num = 32'b00000000001111111111110000000000;
            3:drom_data_num = 32'b00000000111111111111111100000000;
            4:drom_data_num = 32'b00000001111111111111111110000000;
            5:drom_data_num = 32'b00000011111111111111111111000000;
            6:drom_data_num = 32'b00000111111111111111111111100000;
            7:drom_data_num = 32'b00001111111111111111111111110000;
            8:drom_data_num = 32'b00011111111111111111111111111000;
            9:drom_data_num = 32'b00011111111111111111111111111000;
           10:drom_data_num = 32'b00111111111111111111111111111100;
           11:drom_data_num = 32'b00111111111111111111111111111100;
           12:drom_data_num = 32'b00111111111111111111111111111100;
           13:drom_data_num = 32'b01111111111111111111111111111110;
           14:drom_data_num = 32'b01111111111111111111111111111110;
           15:drom_data_num = 32'b01111111111111111111111111111110;
           16:drom_data_num = 32'b01111111111111111111111111111110;
           17:drom_data_num = 32'b01111111111111111111111111111110;
           18:drom_data_num = 32'b01111111111111111111111111111110;
           19:drom_data_num = 32'b00111111111111111111111111111100;
           20:drom_data_num = 32'b00111111111111111111111111111100;
           21:drom_data_num = 32'b00111111111111111111111111111100;
           22:drom_data_num = 32'b00011111111111111111111111111000;
           23:drom_data_num = 32'b00011111111111111111111111111000;
           24:drom_data_num = 32'b00001111111111111111111111110000;
           25:drom_data_num = 32'b00000111111111111111111111100000;
           26:drom_data_num = 32'b00000011111111111111111111000000;
           27:drom_data_num = 32'b00000001111111111111111110000000;
           28:drom_data_num = 32'b00000000111111111111111100000000;
           29:drom_data_num = 32'b00000000001111111111110000000000;
           30:drom_data_num = 32'b00000000000001111110000000000000;
           31:drom_data_num = 32'b00000000000000000000000000000000;
        endcase
 end
 
 endmodule