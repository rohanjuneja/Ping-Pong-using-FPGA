`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 23.10.2016 13:28:25
// Design Name: 
// Module Name: font_player1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module word_player1(
    input [4:0] drom_addr_num,
    output reg [0:223] drom_data_num
);

always @(*)
  begin 
    case (drom_addr_num)
       0:drom_data_num = 224'b01111111111111111111111111110000010000000000000000000000000000000000011111111111111111111110000001000000000000000000000000000010000001111111111111111111111111100111111111111111111111111111000000000000000000000000000000000010;
       1:drom_data_num = 224'b01000000000000000000000000001000010000000000000000000000000000000001000000000000000000000000100001000000000000000000000000000010000010000000000000000000000000000100000000000000000000000000100000000000000000000000000000000110;
       2:drom_data_num = 224'b01000000000000000000000000000100010000000000000000000000000000000010000000000000000000000000010001000000000000000000000000000010000100000000000000000000000000000100000000000000000000000000010000000000000000000000000000001010;
       3:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000010010;
       4:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000100010;
       5:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000001000010;
       6:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000010000010;
       7:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000100000010;
       8:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000001000000010;
       9:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000010000000010;
      10:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      11:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      12:drom_data_num = 224'b01000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001001000000000000000000000000000010010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      13:drom_data_num = 224'b01000000000000000000000000000100010000000000000000000000000000000100000000000000000000000000001000100000000000000000000000000100001000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000010;
      14:drom_data_num = 224'b01000000000000000000000000001000010000000000000000000000000000000100000000000000000000000000001000010000000000000000000000001000000100000000000000000000000000000100000000000000000000000000100000000000000000000000000000000010;
      15:drom_data_num = 224'b01111111111111111111111111110000010000000000000000000000000000000111111111111111111111111111111000000111111111111111111111100000000001111111111111111111111111100111111111111111111111111111000000000000000000000000000000000010;
      16:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000000100000000000000000000000000000100000000000000000000100000000000000000000000000000000000000010;
      17:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000001000000000000000000000000000000100000000000000000000010000000000000000000000000000000000000010;
      18:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000001000000000000000000000000000000000000010;
      19:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000100000000000000000000000000000000000010;
      20:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000010000000000000000000000000000000000010;
      21:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000001000000000000000000000000000000000010;
      22:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000000100000000000000000000000000000000010;
      23:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000000010000000000000000000000000000000010;
      24:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      25:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      26:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      27:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      28:drom_data_num = 224'b01000000000000000000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000010000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      29:drom_data_num = 224'b01000000000000000000000000000000001000000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000001000000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      30:drom_data_num = 224'b01000000000000000000000000000000000100000000000000000000000000000100000000000000000000000000001000000000000000001000000000000000000100000000000000000000000000000100000000000000000000000000001000000000000000000000000000000010;
      31:drom_data_num = 224'b01000000000000000000000000000000000001111111111111111111111111100100000000000000000000000000001000000000000000001000000000000000000001111111111111111111111111100100000000000000000000000000001000000000000000000000000000000010;
    endcase
  end

endmodule