`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/19/2016 06:24:17 PM
// Design Name: 
// Module Name: font_number
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module font_number(
    input [3:0] num_ip,
    input [4:0] drom_addr_num,
    output reg [0:31] drom_data_num
    );
    
always @(*)
    begin
        if(num_ip==4'd0)
        begin
        case (drom_addr_num)
            0:drom_data_num = 32'b00000011111111111111111111000000;
            1:drom_data_num = 32'b00000100000000000000000000100000;
            2:drom_data_num = 32'b00001000000000000000000000010000;
            3:drom_data_num = 32'b00010000000000000000000000001000;
            4:drom_data_num = 32'b00100000000000000000000000000100;
            5:drom_data_num = 32'b01000000000000000000000000000010;
            6:drom_data_num = 32'b01000000000000000000000000000010;
            7:drom_data_num = 32'b01000000000000000000000000000010;
            8:drom_data_num = 32'b01000000000000000000000000000010;
            9:drom_data_num = 32'b01000000000000000000000000000010;
           10:drom_data_num = 32'b01000000000000000000000000000010;
           11:drom_data_num = 32'b01000000000000000000000000000010;
           12:drom_data_num = 32'b01000000000000000000000000000010;
           13:drom_data_num = 32'b01000000000000000000000000000010;
           14:drom_data_num = 32'b01000000000000000000000000000010;
           15:drom_data_num = 32'b01000000000000000000000000000010;
           16:drom_data_num = 32'b01000000000000000000000000000010;
           17:drom_data_num = 32'b01000000000000000000000000000010;
           18:drom_data_num = 32'b01000000000000000000000000000010;
           19:drom_data_num = 32'b01000000000000000000000000000010;
           20:drom_data_num = 32'b01000000000000000000000000000010;
           21:drom_data_num = 32'b01000000000000000000000000000010;
           22:drom_data_num = 32'b01000000000000000000000000000010;
           23:drom_data_num = 32'b01000000000000000000000000000010;
           24:drom_data_num = 32'b01000000000000000000000000000010;
           25:drom_data_num = 32'b01000000000000000000000000000010;
           26:drom_data_num = 32'b01000000000000000000000000000010;
           27:drom_data_num = 32'b00100000000000000000000000000100;
           28:drom_data_num = 32'b00010000000000000000000000001000;
           29:drom_data_num = 32'b00001000000000000000000000010000;
           30:drom_data_num = 32'b00000100000000000000000000100000;
           31:drom_data_num = 32'b00000011111111111111111111000000;
        endcase
        end
        
        else if(num_ip==4'd1)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b00000000000000000000000000000010;
             1:drom_data_num = 32'b00000000000000000000000000000110;
             2:drom_data_num = 32'b00000000000000000000000000001010;
             3:drom_data_num = 32'b00000000000000000000000000010010;
             4:drom_data_num = 32'b00000000000000000000000000100010;
             5:drom_data_num = 32'b00000000000000000000000001000010;
             6:drom_data_num = 32'b00000000000000000000000010000010;
             7:drom_data_num = 32'b00000000000000000000000100000010;
             8:drom_data_num = 32'b00000000000000000000001000000010;
             9:drom_data_num = 32'b00000000000000000000010000000010;
            10:drom_data_num = 32'b00000000000000000000000000000010;
            11:drom_data_num = 32'b00000000000000000000000000000010;
            12:drom_data_num = 32'b00000000000000000000000000000010;
            13:drom_data_num = 32'b00000000000000000000000000000010;
            14:drom_data_num = 32'b00000000000000000000000000000010;
            15:drom_data_num = 32'b00000000000000000000000000000010;
            16:drom_data_num = 32'b00000000000000000000000000000010;
            17:drom_data_num = 32'b00000000000000000000000000000010;
            18:drom_data_num = 32'b00000000000000000000000000000010;
            19:drom_data_num = 32'b00000000000000000000000000000010;
            20:drom_data_num = 32'b00000000000000000000000000000010;
            21:drom_data_num = 32'b00000000000000000000000000000010;
            22:drom_data_num = 32'b00000000000000000000000000000010;
            23:drom_data_num = 32'b00000000000000000000000000000010;
            24:drom_data_num = 32'b00000000000000000000000000000010;
            25:drom_data_num = 32'b00000000000000000000000000000010;
            26:drom_data_num = 32'b00000000000000000000000000000010;
            27:drom_data_num = 32'b00000000000000000000000000000010;
            28:drom_data_num = 32'b00000000000000000000000000000010;
            29:drom_data_num = 32'b00000000000000000000000000000010;
            30:drom_data_num = 32'b00000000000000000000000000000010;
            31:drom_data_num = 32'b00000000000000000000000000000010;
        endcase
        end
        
        else if(num_ip==4'd2)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b01111111111111111111111111111100;
             1:drom_data_num = 32'b00000000000000000000000000000010;
             2:drom_data_num = 32'b00000000000000000000000000000010;
             3:drom_data_num = 32'b00000000000000000000000000000010;
             4:drom_data_num = 32'b00000000000000000000000000000010;
             5:drom_data_num = 32'b00000000000000000000000000000010;
             6:drom_data_num = 32'b00000000000000000000000000000010;
             7:drom_data_num = 32'b00000000000000000000000000000010;
             8:drom_data_num = 32'b00000000000000000000000000000010;
             9:drom_data_num = 32'b00000000000000000000000000000010;
            10:drom_data_num = 32'b00000000000000000000000000000010;
            11:drom_data_num = 32'b00000000000000000000000000000010;
            12:drom_data_num = 32'b00000000000000000000000000000010;
            13:drom_data_num = 32'b00000000000000000000000000000010;
            14:drom_data_num = 32'b00000000000000000000000000000010;
            15:drom_data_num = 32'b00111111111111111111111111111100;
            16:drom_data_num = 32'b01000000000000000000000000000000;
            17:drom_data_num = 32'b01000000000000000000000000000000;
            18:drom_data_num = 32'b01000000000000000000000000000000;
            19:drom_data_num = 32'b01000000000000000000000000000000;
            20:drom_data_num = 32'b01000000000000000000000000000000;
            21:drom_data_num = 32'b01000000000000000000000000000000;
            22:drom_data_num = 32'b01000000000000000000000000000000;
            23:drom_data_num = 32'b01000000000000000000000000000000;
            24:drom_data_num = 32'b01000000000000000000000000000000;
            25:drom_data_num = 32'b01000000000000000000000000000000;
            26:drom_data_num = 32'b01000000000000000000000000000000;
            27:drom_data_num = 32'b01000000000000000000000000000000;
            28:drom_data_num = 32'b01000000000000000000000000000000;
            29:drom_data_num = 32'b01000000000000000000000000000000;
            30:drom_data_num = 32'b01000000000000000000000000000000;
            31:drom_data_num = 32'b00111111111111111111111111111100;
        endcase
        end

        else if(num_ip==4'd3)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b01111111111111111111111111111100;
             1:drom_data_num = 32'b00000000000000000000000000000010;
             2:drom_data_num = 32'b00000000000000000000000000000010;
             3:drom_data_num = 32'b00000000000000000000000000000010;
             4:drom_data_num = 32'b00000000000000000000000000000010;
             5:drom_data_num = 32'b00000000000000000000000000000010;
             6:drom_data_num = 32'b00000000000000000000000000000010;
             7:drom_data_num = 32'b00000000000000000000000000000010;
             8:drom_data_num = 32'b00000000000000000000000000000010;
             9:drom_data_num = 32'b00000000000000000000000000000010;
            10:drom_data_num = 32'b00000000000000000000000000000010;
            11:drom_data_num = 32'b00000000000000000000000000000010;
            12:drom_data_num = 32'b00000000000000000000000000000010;
            13:drom_data_num = 32'b00000000000000000000000000000010;
            14:drom_data_num = 32'b00000000000000000000000000000010;
            15:drom_data_num = 32'b01111111111111111111111111111100;
            16:drom_data_num = 32'b00000000000000000000000000000010;
            17:drom_data_num = 32'b00000000000000000000000000000010;
            18:drom_data_num = 32'b00000000000000000000000000000010;
            19:drom_data_num = 32'b00000000000000000000000000000010;
            20:drom_data_num = 32'b00000000000000000000000000000010;
            21:drom_data_num = 32'b00000000000000000000000000000010;
            22:drom_data_num = 32'b00000000000000000000000000000010;
            23:drom_data_num = 32'b00000000000000000000000000000010;
            24:drom_data_num = 32'b00000000000000000000000000000010;
            25:drom_data_num = 32'b00000000000000000000000000000010;
            26:drom_data_num = 32'b00000000000000000000000000000010;
            27:drom_data_num = 32'b00000000000000000000000000000010;
            28:drom_data_num = 32'b00000000000000000000000000000010;
            29:drom_data_num = 32'b00000000000000000000000000000010;
            30:drom_data_num = 32'b00000000000000000000000000000010;
            31:drom_data_num = 32'b01111111111111111111111111111100;
        endcase
        end
        
        else if(num_ip==4'd4)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b01000000000000000000000000000010;
             1:drom_data_num = 32'b01000000000000000000000000000010;
             2:drom_data_num = 32'b01000000000000000000000000000010;
             3:drom_data_num = 32'b01000000000000000000000000000010;
             4:drom_data_num = 32'b01000000000000000000000000000010;
             5:drom_data_num = 32'b01000000000000000000000000000010;
             6:drom_data_num = 32'b01000000000000000000000000000010;
             7:drom_data_num = 32'b01000000000000000000000000000010;
             8:drom_data_num = 32'b01000000000000000000000000000010;
             9:drom_data_num = 32'b01000000000000000000000000000010;
            10:drom_data_num = 32'b01000000000000000000000000000010;
            11:drom_data_num = 32'b01000000000000000000000000000010;
            12:drom_data_num = 32'b01000000000000000000000000000010;
            13:drom_data_num = 32'b01000000000000000000000000000010;
            14:drom_data_num = 32'b01000000000000000000000000000010;
            15:drom_data_num = 32'b00111111111111111111111111111100;
            16:drom_data_num = 32'b00000000000000000000000000000010;
            17:drom_data_num = 32'b00000000000000000000000000000010;
            18:drom_data_num = 32'b00000000000000000000000000000010;
            19:drom_data_num = 32'b00000000000000000000000000000010;
            20:drom_data_num = 32'b00000000000000000000000000000010;
            21:drom_data_num = 32'b00000000000000000000000000000010;
            22:drom_data_num = 32'b00000000000000000000000000000010;
            23:drom_data_num = 32'b00000000000000000000000000000010;
            24:drom_data_num = 32'b00000000000000000000000000000010;
            25:drom_data_num = 32'b00000000000000000000000000000010;
            26:drom_data_num = 32'b00000000000000000000000000000010;
            27:drom_data_num = 32'b00000000000000000000000000000010;
            28:drom_data_num = 32'b00000000000000000000000000000010;
            29:drom_data_num = 32'b00000000000000000000000000000010;
            30:drom_data_num = 32'b00000000000000000000000000000010;
            31:drom_data_num = 32'b00000000000000000000000000000010;
        endcase
        end
            
        else if(num_ip==4'd5)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b00111111111111111111111111111110;
             1:drom_data_num = 32'b01000000000000000000000000000000;
             2:drom_data_num = 32'b01000000000000000000000000000000;
             3:drom_data_num = 32'b01000000000000000000000000000000;
             4:drom_data_num = 32'b01000000000000000000000000000000;
             5:drom_data_num = 32'b01000000000000000000000000000000;
             6:drom_data_num = 32'b01000000000000000000000000000000;
             7:drom_data_num = 32'b01000000000000000000000000000000;
             8:drom_data_num = 32'b01000000000000000000000000000000;
             9:drom_data_num = 32'b01000000000000000000000000000000;
            10:drom_data_num = 32'b01000000000000000000000000000000;
            11:drom_data_num = 32'b01000000000000000000000000000000;
            12:drom_data_num = 32'b01000000000000000000000000000000;
            13:drom_data_num = 32'b01000000000000000000000000000000;
            14:drom_data_num = 32'b01000000000000000000000000000000;
            15:drom_data_num = 32'b00111111111111111111111111111100;
            16:drom_data_num = 32'b00000000000000000000000000000010;
            17:drom_data_num = 32'b00000000000000000000000000000010;
            18:drom_data_num = 32'b00000000000000000000000000000010;
            19:drom_data_num = 32'b00000000000000000000000000000010;
            20:drom_data_num = 32'b00000000000000000000000000000010;
            21:drom_data_num = 32'b00000000000000000000000000000010;
            22:drom_data_num = 32'b00000000000000000000000000000010;
            23:drom_data_num = 32'b00000000000000000000000000000010;
            24:drom_data_num = 32'b00000000000000000000000000000010;
            25:drom_data_num = 32'b00000000000000000000000000000010;
            26:drom_data_num = 32'b00000000000000000000000000000010;
            27:drom_data_num = 32'b00000000000000000000000000000010;
            28:drom_data_num = 32'b00000000000000000000000000000010;
            29:drom_data_num = 32'b00000000000000000000000000000010;
            30:drom_data_num = 32'b00000000000000000000000000000010;
            31:drom_data_num = 32'b01111111111111111111111111111100;
        endcase
        end
            
        else if(num_ip==4'd6)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b00111111111111111111111111111100;
             1:drom_data_num = 32'b01000000000000000000000000000000;
             2:drom_data_num = 32'b01000000000000000000000000000000;
             3:drom_data_num = 32'b01000000000000000000000000000000;
             4:drom_data_num = 32'b01000000000000000000000000000000;
             5:drom_data_num = 32'b01000000000000000000000000000000;
             6:drom_data_num = 32'b01000000000000000000000000000000;
             7:drom_data_num = 32'b01000000000000000000000000000000;
             8:drom_data_num = 32'b01000000000000000000000000000000;
             9:drom_data_num = 32'b01000000000000000000000000000000;
            10:drom_data_num = 32'b01000000000000000000000000000000;
            11:drom_data_num = 32'b01000000000000000000000000000000;
            12:drom_data_num = 32'b01000000000000000000000000000000;
            13:drom_data_num = 32'b01000000000000000000000000000000;
            14:drom_data_num = 32'b01000000000000000000000000000000;
            15:drom_data_num = 32'b00111111111111111111111111111100;
            16:drom_data_num = 32'b01000000000000000000000000000010;
            17:drom_data_num = 32'b01000000000000000000000000000010;
            18:drom_data_num = 32'b01000000000000000000000000000010;
            19:drom_data_num = 32'b01000000000000000000000000000010;
            20:drom_data_num = 32'b01000000000000000000000000000010;
            21:drom_data_num = 32'b01000000000000000000000000000010;
            22:drom_data_num = 32'b01000000000000000000000000000010;
            23:drom_data_num = 32'b01000000000000000000000000000010;
            24:drom_data_num = 32'b01000000000000000000000000000010;
            25:drom_data_num = 32'b01000000000000000000000000000010;
            26:drom_data_num = 32'b01000000000000000000000000000010;
            27:drom_data_num = 32'b01000000000000000000000000000010;
            28:drom_data_num = 32'b01000000000000000000000000000010;
            29:drom_data_num = 32'b01000000000000000000000000000010;
            30:drom_data_num = 32'b01000000000000000000000000000010;
            31:drom_data_num = 32'b00111111111111111111111111111100;
        endcase
        end
            
        else if(num_ip==4'd7)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b01111111111111111111111111111100;
             1:drom_data_num = 32'b00000000000000000000000000000010;
             2:drom_data_num = 32'b00000000000000000000000000000010;
             3:drom_data_num = 32'b00000000000000000000000000000010;
             4:drom_data_num = 32'b00000000000000000000000000000010;
             5:drom_data_num = 32'b00000000000000000000000000000010;
             6:drom_data_num = 32'b00000000000000000000000000000010;
             7:drom_data_num = 32'b00000000000000000000000000000010;
             8:drom_data_num = 32'b00000000000000000000000000000010;
             9:drom_data_num = 32'b00000000000000000000000000000010;
            10:drom_data_num = 32'b00000000000000000000000000000010;
            11:drom_data_num = 32'b00000000000000000000000000000010;
            12:drom_data_num = 32'b00000000000000000000000000000010;
            13:drom_data_num = 32'b00000000000000000000000000000010;
            14:drom_data_num = 32'b00000000000000000000000000000010;
            15:drom_data_num = 32'b00000000000000000000000000000010;
            16:drom_data_num = 32'b00000000000000000000000000000010;
            17:drom_data_num = 32'b00000000000000000000000000000010;
            18:drom_data_num = 32'b00000000000000000000000000000010;
            19:drom_data_num = 32'b00000000000000000000000000000010;
            20:drom_data_num = 32'b00000000000000000000000000000010;
            21:drom_data_num = 32'b00000000000000000000000000000010;
            22:drom_data_num = 32'b00000000000000000000000000000010;
            23:drom_data_num = 32'b00000000000000000000000000000010;
            24:drom_data_num = 32'b00000000000000000000000000000010;
            25:drom_data_num = 32'b00000000000000000000000000000010;
            26:drom_data_num = 32'b00000000000000000000000000000010;
            27:drom_data_num = 32'b00000000000000000000000000000010;
            28:drom_data_num = 32'b00000000000000000000000000000010;
            29:drom_data_num = 32'b00000000000000000000000000000010;
            30:drom_data_num = 32'b00000000000000000000000000000010;
            31:drom_data_num = 32'b00000000000000000000000000000010;
        endcase
        end
        
        else if(num_ip==4'd8)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b00111111111111111111111111111100;
             1:drom_data_num = 32'b01000000000000000000000000000010;
             2:drom_data_num = 32'b01000000000000000000000000000010;
             3:drom_data_num = 32'b01000000000000000000000000000010;
             4:drom_data_num = 32'b01000000000000000000000000000010;
             5:drom_data_num = 32'b01000000000000000000000000000010;
             6:drom_data_num = 32'b01000000000000000000000000000010;
             7:drom_data_num = 32'b01000000000000000000000000000010;
             8:drom_data_num = 32'b01000000000000000000000000000010;
             9:drom_data_num = 32'b01000000000000000000000000000010;
            10:drom_data_num = 32'b01000000000000000000000000000010;
            11:drom_data_num = 32'b01000000000000000000000000000010;
            12:drom_data_num = 32'b01000000000000000000000000000010;
            13:drom_data_num = 32'b01000000000000000000000000000010;
            14:drom_data_num = 32'b01000000000000000000000000000010;
            15:drom_data_num = 32'b00111111111111111111111111111100;
            16:drom_data_num = 32'b01000000000000000000000000000010;
            17:drom_data_num = 32'b01000000000000000000000000000010;
            18:drom_data_num = 32'b01000000000000000000000000000010;
            19:drom_data_num = 32'b01000000000000000000000000000010;
            20:drom_data_num = 32'b01000000000000000000000000000010;
            21:drom_data_num = 32'b01000000000000000000000000000010;
            22:drom_data_num = 32'b01000000000000000000000000000010;
            23:drom_data_num = 32'b01000000000000000000000000000010;
            24:drom_data_num = 32'b01000000000000000000000000000010;
            25:drom_data_num = 32'b01000000000000000000000000000010;
            26:drom_data_num = 32'b01000000000000000000000000000010;
            27:drom_data_num = 32'b01000000000000000000000000000010;
            28:drom_data_num = 32'b01000000000000000000000000000010;
            29:drom_data_num = 32'b01000000000000000000000000000010;
            30:drom_data_num = 32'b01000000000000000000000000000010;
            31:drom_data_num = 32'b00111111111111111111111111111100;
        endcase
        end
        
        else if(num_ip==4'd9)
        begin
        case (drom_addr_num)
             0:drom_data_num = 32'b00111111111111111111111111111100;
             1:drom_data_num = 32'b01000000000000000000000000000010;
             2:drom_data_num = 32'b01000000000000000000000000000010;
             3:drom_data_num = 32'b01000000000000000000000000000010;
             4:drom_data_num = 32'b01000000000000000000000000000010;
             5:drom_data_num = 32'b01000000000000000000000000000010;
             6:drom_data_num = 32'b01000000000000000000000000000010;
             7:drom_data_num = 32'b01000000000000000000000000000010;
             8:drom_data_num = 32'b01000000000000000000000000000010;
             9:drom_data_num = 32'b01000000000000000000000000000010;
            10:drom_data_num = 32'b01000000000000000000000000000010;
            11:drom_data_num = 32'b01000000000000000000000000000010;
            12:drom_data_num = 32'b01000000000000000000000000000010;
            13:drom_data_num = 32'b01000000000000000000000000000010;
            14:drom_data_num = 32'b01000000000000000000000000000010;
            15:drom_data_num = 32'b00111111111111111111111111111100;
            16:drom_data_num = 32'b00000000000000000000000000000010;
            17:drom_data_num = 32'b00000000000000000000000000000010;
            18:drom_data_num = 32'b00000000000000000000000000000010;
            19:drom_data_num = 32'b00000000000000000000000000000010;
            20:drom_data_num = 32'b00000000000000000000000000000010;
            21:drom_data_num = 32'b00000000000000000000000000000010;
            22:drom_data_num = 32'b00000000000000000000000000000010;
            23:drom_data_num = 32'b00000000000000000000000000000010;
            24:drom_data_num = 32'b00000000000000000000000000000010;
            25:drom_data_num = 32'b00000000000000000000000000000010;
            26:drom_data_num = 32'b00000000000000000000000000000010;
            27:drom_data_num = 32'b00000000000000000000000000000010;
            28:drom_data_num = 32'b00000000000000000000000000000010;
            29:drom_data_num = 32'b00000000000000000000000000000010;
            30:drom_data_num = 32'b00000000000000000000000000000010;
            31:drom_data_num = 32'b01111111111111111111111111111100;
        endcase
        end
     end
endmodule